	rand bit [2:0]a;
	constraint b_size{a<3;}	//constraint identifiers are different,so no-overriding takes place
endclass

parent p1_h;
child1 ch1_h;

module parent_child_same_prop;

	initial
		begin
			ch1_h = new();

			for(int i=0;i<7;i++)
				begin
					assert(ch1_h.randomize());
					$display("ch1_h: %p",ch1_h);
				end
		end
endmodule


/* output

ch1_h: '{a:'h1, a:'h2}
ch1_h: '{a:'h2, a:'h0}
ch1_h: '{a:'h1, a:'h1}
ch1_h: '{a:'h2, a:'h1}
ch1_h: '{a:'h2, a:'h1}
ch1_h: '{a:'h2, a:'h1}
ch1_h: '{a:'h1, a:'h2}

*/
